�}P8 �'  6z-Fn��Q��� ^:���`<�y��bjneFN�Ƙw��D���1�,��r80��̄��)������ӳ�kUomOD4r��4��s���H�"�T#	0 AUF���J1�-رʹ��eyn>l_�{m'(�'}���mO�I��68RZn	�Prg���V�w񃋂Fcm�#8� c��n��ſ�P�,��gV��A��z&���;���J��q�%��y�VY^���i
�s��fD{�r��ud�+�nݲ;͠ط���G�_8.-�e1)ջ�����'r+�� eZ���So��\��-����a_:�]軠μ��f߆d�ՃY��� :�.�jl��:�TK�FY�{,>٣�'�p�@�L��#�:*
)��ɀdR��p<@�g�K��n��c�QܛVs�/],XX��D�}_��ê���'�s�G8�Z.��:�.s�}�1%����5͗k��d�����n(����"�^p߶ћlDi掌>9���=�M�3�\UN��h��d����N�*�5W�`g����F��P�Ē������a^Z��N�%qf�X�T�1�K,Тgm��Q(#�H��oW��+�i���"r�����("�w�T��pj
#(:l�pmW��^r����D�/*GK�͠�!M'��HR�!( C>[�%�����'L�+����P� 90�9}[�~&�X#֞]I�I�F��R �w�@�􃈲l�n[+�0���f��睨�XQ1��$�a!�2O��cK8&���2z���>(�7�f{���v^��\��3�L���U�gM�-Z�A��H`�p#^e�k��VH����?�7�=�I�owg07�\�6�*�ό2r��|K�em����Х�L�P����į^,�����6�GB���J�8���mT�.��ݩ�B�1~M+��N,��c�5�O�u��L$���x5Q��~�1���LTT�o@iq�Vyɗ&4��-l�"@D��Ӄ`�	[��t��Lk�a��g~e¿�vp|�Vxփ���$�ӨN�o@T�b��jhy�\%1a��2�D_}�Ǟ����Ü�y�Y7��r��O�J�d�`�����/��xZ�g5f�����ə�0��F||��d-@�,�������ִ�_L��lv��ŴJ�_�Y$��g`���>�BS���X��j�@� 1�P�PXí�I�l�^.Ge����p��[��s�u�d�D�N	S���q�
��B��L�],�m��\?B݁�PY��#ȕ�ق�AB ���i�E�gV�h'^�aA�S�g%�U7)��v1�:�r.DuyfR"I"��F�a@x����^76#D�Psw�7Wf���ϛ�8�Q��ń!�BseY?'��j�n��Z��Pɡճ���o�6����l%�'�����7WS����FZ(��O��A�Aɑ�"7�����8�=L}t���e^¢�
�9����J���J��{���]�v�e2s)T�!N[l]/<��C��d���
��
��6�3�6��ܡ��ܶV!�
�o��ޟ�
QIwb'���X���
51�RV��@�����V���u쥩`K�6	OCQ7�hD���3�`t�F����ԩ���[���VNIs�OLӽ�_Kd����ӏ��gC	`Yc��k�*ܵ)�������0�)b�����?�^p�ǭ0}�x���퉾�Ě�`��%���3s�M��Ĕ�1�d�f����0�='?Ų?႔��<�C�-��F%�W�+�MK������K�V�%���@T��zv�.�B��`W��җuz$7���*�����~�A�zF�����g�l���7%��r�����L���U�Vs��xFJ�[����~
�OʸY�����8��HO�h#X�|3"�خ)_G��(5�jދ��1��� ~�[��3�Uc��ό�$h��1�\��D��k3@[ӔC8�#3�j�ʷmޏt �6c�ڒH��\�q�l�:g<r�-~R�}�p��^�3-4��ɠN��P��:���@���08��R~ҁw�Y����	'Pr y��U�"E��1�Ϗ������z�f����P���Aqelx;+[���S'(W2�g�PNr�]6�z��EN!d��֓o�5�����q�0ٓϸ�W��x�L�6�w�-�E���Q�9]\���,��cS2X ��p�R�SXJ��Q��:it�
A1�^JBؤ��N`u��Л�otX�Ȍj私>����z8�LwS�����+���~W�M���y�o�����b�1s/���	�Y#��,>��^U�U��d�jɜU��N� 5	�|I�7.Kr)�7�X�z�s��Z�]���ʵ�����3N}���W���a^''�yS�$Ɗ8�D��Sp��ߋp)Y��dW�m.�G�
�&�*�0˹3�eO�h�9k����#���5��gef�Yr��vU������~�>�6)�C�
�C>7�8X���|���q�(Զ'�Kxl '4�	�<(,��M����\�~�ԦB���׸R��&��{���!��t-G���rA"���"����%V�Lu��m2&|����BN�ӖC��p�i�U��d"'��) o�Q~Q;�"b��[x���u��*����rs��zt��vL_��'�A)��SǏm?��+��;b�� ���6���t\����< -g�܄�tF�F��Ĵ,��Ubj�P�$�E�9����
�L�Wa��ôZ���#���%hh�����{F�$sES��1@A���<�ƥfnLO��t�$��>	і�K���r	а)��%�Kl�D�8�����(-"�
����=��hl�-��7)�BPih�$�HP<_�9q�/��f�Z5�fևq��Z���u���qx,��C��q/[�1�k:o��Z�ת��YQέ��XF�Gi�#�U����į������9Bb?--d*wK�ҥ+d��6��7l�����_fFIO��5��=��Ǐ/=�ޜ��4�l]/<]����=fxI������"vG�
9�[T'`(Ñ8h�g��!�ɱ�PbP;9�����b�W�l����!MR�MA�zWE��*����c|�S�~s��`�oF��F����Ԙ���i������h��A�ϖ�C�Þ嶗n[rD /��k�*ܵ)�������*�x�f��s�Q��s!��R7�������d���`�|(���'w�I�+��~���L�%�sDE�͒�'�&%xd_��f�����Y�,�T��}"L�2�&�@\�j�Ô&�f�����m���`s��"/�v�f��D?s3����Q:V{�ض�s�ؤ��^�e�"�����C� H�����<�5����M�Ӏ9�Qm��RFlU?_��N3�n�"A:�������=G����o�(�R�Pi��
�;NZ����*e,�����F�\4�1G�V�ezM��ܑeX��@U�,�y�jÌp4�6 K_��ν�|u�X����t�ip�GuZ���l#��:���&����aP���/�1l�zG*��}#�t]��Ǔ4��vE����t��ل�\�hٓ��ݦ�ؐ��
ީ�KЉۋ��i�"�Z�~��oG�n��>�!�z���w�M��o�ԁ`(�ŶFCj��o�}��.Q�Vr�{Ex�!���z��b��[3J�|����M4�ꤴ�I��~}XO�sk\��4��d}Wr@a6"u6�o2��w��f����i@�(�4aS��-^V�@�x��>}��D�i�0�ɓ�.�\�&D��bd�b�y2�"��${�8�5��D��hX��SN��)05��S�v�Z�=/-͝}��ߴѺJl������ �����;�}�|���VT�%
�-�5�.I$q��=�D$ G>��{�N��̞�'���+���,ɤ]���k�^��s��RF%ʄ��� 㻨��B�VY�Ъ�����s�����X$ĉw�a��eO�H�n�m?T�r�Z��^��`=�rxBlD���(����P���;��\K�����f9�GZ,�"�L����0��M�I-v��Ec�9Dx(;�
��'z��\�`ڢzp�>݅�1#����#������ϛ%�<
�m����֍@�{�f�a�B�&�Q@n��>�j�θ�M�� iV]y-�@�`	�����<?��a�>��[ �Y!}�W�p�ʩԤ#\���S&�}ł�y�aא��
�Qh�\�ҚFN�'����uX�5y��f]twD�����0Q��Z����=&K/m*K��;���;�A��+��t̘e8[q�����[�o�'�}�AB�:XE[�Q��"�*��2赡u��N��\���b��n=ΒfB�Eh�@�C���0�C�f�����"�V4�̀??�b�2�~Us��4�@�=�$~�,���6!�8���I�NY�
K��<�wW҉�us��v�d�����ˁ��|��冻��e{�2^E#M�uN=�**~dM�ֱ4�d&s�����l#��:-�%";�!�#bG��׼�"U��s����!�w����z����7jz�T�n�.d�r�!@3G��9-'��"��� +P��2Gˍ���{'�DM8M���V�(4����2R��+�"�=e��9£��ߡ�o�}��xG&�l_�	0�~h���H��b�^LK�{����E#R^���68�q�{�Z}`�2fM��u��,/p}Zt	>*YH�v%)��^��`����.�[�y!SW�}�F@�W�U�$:��D��8��4�g�#	3��BDD�1�7w�ګ�T���=��:��;*��#99�O�uO�)��9�U���˘�Dʦ"��&�ځr�U����+�t�U#��A�=/�s�b�e�#^)'��s�rs|��j@����;�'�1f�'��P0�h���h�)�/�􉀖�#��:��	[{�#�e/�4J�f䒕A	Ebq�q*�=��� և��4}��]/ �M��&�����bs��	�P�hlD$9�	hn�� ����v.R?sMn��Y������Q)��ɦj�zA�Z?%���f�j�OR_���)���+�y�?)�7�A(����M���-�?岿a���/�U��ߟ��o�Q֭�"@e|�����I
E=-����p�
���E�/ ��܀����J��Ǭ�GK���0����\SY��O��7E̚�aK���z4N{�^�
��7�c�l��q�V�����������A���UgI��2��	x}�م$����&Qn�A�,vIW�>�Ý�փ����'{a]��HT�`d��V �].V_D���"�Ip�%h����aKp�Q���`�Y���S*�A��8�:�����{>�Cq�=�ZiAS��x_��3l_L��z����j��V�}�'ER,B�XW��C%Q���ͨ	Gw�FګiL��Hkd��@.��7 ˡ�z�+~��/��em!���6Pa���F�!br���I|����^�u�c�lD*|`�4�g�	��?܂7�cX�O�,-��jǛ��η��4�[�^�B7B���򏾅�y�K���l�d��A�f�:�3�ރ��AS�x�t��[���'�%l�8�sVӬ��T'W0�C�E7���S�xy�/�	�5�aZ�tX�i�uGƣ���\^`.^�߇�,}��!�0��-#6�ڱ���Ը��z�����h�Yk�E�+J�*5�O�ߣ��k�\- ���zEv&,E�A�;B����Ӳ���/D =;���I"���	a���u�YDQ&Y6m��GtV�|-)w�D`��^��=�4�n05&zzb��Ռr�~
�⁒��>F��8�X�#_/`�)'x�m�L�Uƌsz����m�2nY^"}mn�= n�l�w�����	ºP�S&$V�%��(�o��q�[ ;Re.�$����k�!U��`�ކ�j�����ER���|�Dܳ�۠��0�ir:8U����'�nB;?�h���NP��"�`%n�vX�L�l�#-��Æ� _�<����bۿ���"`[����� bb�M4��C��CC,
��D�)RarR�n�s�g�r�[��E��ɰϛ5EAm|2�.��#g˔`����.6�;���j���Ƣ2���̴�6�dx6c�G��&�'j9��ȅ˛��'9e�ǰ
^U�%�%����ќk�`��u'�u1���*#7'�"~��;�`DQn@�V!H{(i�
ȹ0 Ū�$J�)��eI��A�!r�u��y�-�g�z�e(�H<&����rO� ��n�����=��[��6��$`�z�(ڑn�l�=�.�e���I�V�?fM�:o}R%��]�_�-O�n#�F�:ܵ8u<?�u��tuՎ�寻&��m��M�)�.|��>����V�0�ԏ�8.tG?f��(�I�R>���t���=�4��/�x*F���?�R>4	T���
�$���ﳴK@y�d������,%���x����A�U��T��N��V�^{���	�S��l�+�A����w�߅�@�2�s̫"B�kĚ�BEAn
�����&�t� +X��w���D
�i��s���7�!". Pf�J��c�X�x�������Y���X�\Tv��j4ސH'K�\�'�?؛>aϯ�ₕ�Dd?d	?�6�<���D�@�` Z01�$���
�S���*%��i?��YG�pL�2��͊����<��� �U��~k������4S�1q;~�� �і7���0��~�邜��%[xм��9�W��R�rԛ�и����,��y���>� ^�5�sDn�7a}����+�ݨ�L@t�E{7^�f�mP7}���P���������Gˠy	8�ڑJg�N��JQ��	y���TS:�]E+ À�V�&�f���~ȇdU~N�������B��0�đ۹|�����	_�P�e��`�-�D^�pP�6Q�z����e�/ڃ��h�f��ؠ/w��dT�HV�g�R3����%�Q�U����!���/l�$�6kr��C;ًZbߖ0NR�Mٴ�7T<6�;���w�]�dÙ�N��DQKTY5?�vA��-�rCK��pܴ�n�u� �4�fL�] {.?��	'{<<�/�*�hQ*�����(K�d����3�R�����M9\��b�:N%��M�m�3��咩w0#c�K�Ⰺ��M��.E���յ�q?���
K.��ZeI ~T�)dS=���ZQ��+�}��U�xf=�`U���4�`W�~	hZģ�����H�L��a3R���R�]���;1��w:1O�!wg��9�e*�C@�km�V3y��:_��rI�������g}&W�Ǩ*UO��R\�[K���{����gʩ�jx���2oL#����y���U6nm����a�"M0�5����_Kc��j��I���P��ߣ�vüm�|�[@&*|ƚ:���Ri�1<�ǧO>���w�[��B>4�t�e���2����g�S�oT3��rҋ��m�X������2�%ʢy΄+l&��P�6D�N�el��P�*�� �E����,���$�HO�	ɩ;��9�)6��j}��*�����Eb��[S�0�.I�]q8B��Uĳ�M��ZI�l�X���n�$�����" J筺���M`օv !��O�6Q=1k��0�.��s?̤����c -�ĺ�HF��?ʼV�dX��'��YXRKn�:�>�E� ;5A��&��F7h���Ò���C��#�y�n.�B6��Y-�9v?4��F�ޔV��L,�hɵ/�'����-�59��}X�l���_�귯�i!�r%]�} h�Q��I�#���q
f���M�� a)2�n�#�nBT��}m���*�f���z&J]���~���ĵ���C�U�m�h�����EfOq�͹O/���[~�Ib&",����H.=��_Y��_!>�����A�8:�m�%RA���vݽV<]�F�K�KkJJ�ا/\�>�ֲ�Y�����l�k�r=��?�'�y�W#ّ!��l#��:� ��	m�QZ|�U������ٺW�d���R)/)���.zJ�Y��:d���A8j��8���p�P��T�/M�&���LE=�����C#���>p�>��o�-S�Ȏ�5�����`���Ԅ����i���o�}��uT5�/�{Hd�6���^��F��EA�%ٌ�n�b����e�q�:�6(.�~k@��9��r])4X8/;TS�jZp���m����d\�?� DEw�>Y�_��X��V|7��I�
�J����F�!�kT>���~�n?�R��$�3���U��>��v ��|��2�u�7�N(�8<��睎�/o��q�������*�n���O�I��7H��;�TV�%
�-�5�.I$q��=�D$ G>����:�`��-&�K-����!8�CnE�E�	�P��D�Q��Y����6��䍚�[��6��<Y޺��Tg/6r��8Q�q�&ТI߭#R�ܫuu-kN����p־l�"�����U�uC����p<Rm��FWD4�kn��.�o�
a�o��B U1�QH4������W��]m ���2:�
��_J*���/�.�R�ja1��u�G'����!dV�$m�U�Cr+ �qU��G��__��zc��%�%�D�?W��RI�Ѧ����j�	�6'
ϳՍA�gǞ��e��X^�5�ߋTyY}�z����ʌ}؇�)fG���N�ͬ"b���)����e>J�ʽ�A�+%���뱨(A��cIp�<�^<tV���v�V�!T}�d?��9��>g��R����׈���M��q�a�s�en���A����H�f���m.�&t�E��k��|�_v������_���_}_���]ՠ_��hD�7��	 Vm�9��=���٬��5��Z���Z5��S�Q�P���f��{��W�@�����Q�F��xo�� A��)�t����۫C�P48�pv7�����ۯ����edu�H�ɼ_BYTE_POS_WIDTH{1'b0}};
			r.next_byte_flag	<= 1'b0;
			r.trans_en			<= 1'b0;
			r.first_ofs			<= {CONV_OFS_WIDTH{1'b0}};
		end
	end

endmodule

//--------------------------------------------------------------------------------------------------
// eof
//--------------------------------------------------------------------------------------------------

